package dma_pkg;
  `include "uvm_macros.svh"
	 import uvm_pkg::*;
	`include "dma_sequence_item.sv"
	`include "dma_intr_register.sv"
	`include "dma_ctrl_register.sv"
	`include "dma_io_addr_register.sv"
	`include "dma_mem_addr_register.sv"
	`include "dma_extra_info_register.sv"
	`include "dma_status_register.sv"
	`include "dma_transfer_count_register.sv"
	`include "dma_descriptor_addr_register.sv"
	`include "dma_error_status_register.sv"
	`include "dma_configure_register.sv"
	`include "dma_reg_file.sv"
	`include "dma_reg_block.sv"
	`include "dma_ctrl_sequence.sv"
	`include "dma_regression_sequence.sv"
	`include "dma_report_server.sv"
	`include "dma_adapter.sv"
	`include "dma_sequencer.sv"
	`include "dma_driver.sv"
	`include "dma_monitor.sv"
	`include "dma_agent.sv"
	`include "dma_subscriber.sv"
	`include "dma_environment.sv"
	`include "dma_test.sv"
endpackage

